library verilog;
use verilog.vl_types.all;
entity full_adder_1bit_tb_v is
end full_adder_1bit_tb_v;
