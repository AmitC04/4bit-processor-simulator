library verilog;
use verilog.vl_types.all;
entity alu_4bit_tb_v is
end alu_4bit_tb_v;
