library verilog;
use verilog.vl_types.all;
entity ram_16x4_sync_tb_v is
end ram_16x4_sync_tb_v;
