library verilog;
use verilog.vl_types.all;
entity adder_4bit_tb_v is
end adder_4bit_tb_v;
