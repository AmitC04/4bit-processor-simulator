library verilog;
use verilog.vl_types.all;
entity registered_alu_tb_v is
end registered_alu_tb_v;
