library verilog;
use verilog.vl_types.all;
entity processor_4bit_tb_v is
end processor_4bit_tb_v;
