library verilog;
use verilog.vl_types.all;
entity instruction_decoder_tb_v is
end instruction_decoder_tb_v;
