library verilog;
use verilog.vl_types.all;
entity half_adder_tb_v is
end half_adder_tb_v;
