library verilog;
use verilog.vl_types.all;
entity xor_gate_tb_v is
end xor_gate_tb_v;
