library verilog;
use verilog.vl_types.all;
entity processor_4bit_tb is
end processor_4bit_tb;
